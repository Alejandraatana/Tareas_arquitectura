--Alejandra Rodriguez Sanchez Ing. en Computacion

